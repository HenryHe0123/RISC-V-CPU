//Reservation Station

module RS(

);

endmodule