//Registers

module registers(

);

endmodule