//Instruction Fetcher

module IFetcher(
    input wire clk, rst, rdy
    
);

endmodule