//Register File

module regFile(

);

endmodule