//Load Store Buffer

module LSB(

);

endmodule