//Predictor

module predictor(
    input wire clk, rst, rdy,
    output wire predict
);

assign predict = 1'b1;

endmodule