//Reorder Buffer

module ROB(

);

endmodule