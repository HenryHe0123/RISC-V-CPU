//Memory Controller

module mem_controller(
    
);

endmodule