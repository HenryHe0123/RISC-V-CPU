//Instruction Queue (Issue)

module IQueue(

);

endmodule